module dca_tb;

endmodule