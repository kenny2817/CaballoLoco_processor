import alu_pkg::*;

module alu #(
    parameter DATA_WIDTH
) (
    input logic [DATA_WIDTH - 1 : 0]    i_elemA,
    input logic [DATA_WIDTH - 1 : 0]    i_elemB,
    input alu_op_e                      i_op,
    output logic [DATA_WIDTH - 1 : 0]   o_output
);
    always_comb begin
        case (i_op)
            ADD:        o_output = (i_elemA + i_elemB);
            SUB:        o_output = (i_elemA - i_elemB);
            AND:        o_output = (i_elemA & i_elemB);
             OR:        o_output = (i_elemA | i_elemB);
            XOR:        o_output = (i_elemA ^ i_elemB);
            MUL:        o_output = (i_elemA * i_elemB);
            DIV:        o_output = (i_elemA / i_elemB);
            default:    o_output = 'x;
        endcase
    end
endmodule
