
import cmp_pkg::*;
import alu_pkg::*;
import opcodes_pkg::*;

module cbl



endmodule

module cbl_tb:



endmodule